**.subckt nmos
XM1 vd vg vss vss sky130_fd_pr__nfet_01v8 L='l' W='w' nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult='m' m='m' 
VG vg vss {vg} 
VD vd vss {vdd} 
VSS vss GND {vss} 
**.ends
.GLOBAL GND
** flattened .save nodes
.end
